`include "defines.vh"

module a_register(
    input clk,
    input areset,

    input set,
    input [`WORD_SIZE - 1 : 0] in,
    output [`WORD_SIZE - 1 : 0] out
);
    wire clk;
    wire areset;

    wire set;
    wire [`WORD_SIZE - 1 : 0] in;
    wire [`WORD_SIZE - 1 : 0] out;

    reg [`WORD_SIZE - 1 : 0] a;

    always @(clk) if (set) a <= in;

    assign out = a;
endmodule
